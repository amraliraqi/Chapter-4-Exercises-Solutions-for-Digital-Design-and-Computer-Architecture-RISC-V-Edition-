module ex_14 (
	input [5:0] a,
	output [63:0] y );

     wire [11:0] y2_4;
     ex_13 DU0 (a[1:0], y2_4[3:0]);
     ex_13 DU1 (a[3:2], y2_4[7:4]);
     ex_13 DU2 (a[5:4], y2_4[11:9]);

assign y[0] = y2_4[0] & y2_4[4] & y2_4[8];
assign y[1] = y2_4[1] & y2_4[4] & y2_4[8];
assign y[2] = y2_4[2] & y2_4[4] & y2_4[8];
assign y[3] = y2_4[3] & y2_4[4] & y2_4[8];
assign y[4] = y2_4[0] & y2_4[5] & y2_4[8];
assign y[5] = y2_4[1] & y2_4[5] & y2_4[8];
assign y[6] = y2_4[2] & y2_4[5] & y2_4[8];
assign y[7] = y2_4[3] & y2_4[5] & y2_4[8];

assign y[8] = y2_4[0] & y2_4[6] & y2_4[8];
assign y[9] = y2_4[1] & y2_4[6] & y2_4[8];
assign y[10] = y2_4[2] & y2_4[6] & y2_4[8];
assign y[11] = y2_4[3] & y2_4[6] & y2_4[8];

assign y[12] = y2_4[0] & y2_4[7] & y2_4[8];
assign y[13] = y2_4[1] & y2_4[7] & y2_4[8];
assign y[14] = y2_4[2] & y2_4[7] & y2_4[8];
assign y[15] = y2_4[3] & y2_4[7] & y2_4[8];

assign y[16] = y2_4[0] & y2_4[4] & y2_4[9];
assign y[17] = y2_4[1] & y2_4[4] & y2_4[9];
assign y[18] = y2_4[2] & y2_4[4] & y2_4[9];
assign y[19] = y2_4[3] & y2_4[4] & y2_4[9];

assign y[20] = y2_4[0] & y2_4[5] & y2_4[9];
assign y[21] = y2_4[1] & y2_4[5] & y2_4[9];
assign y[22] = y2_4[2] & y2_4[5] & y2_4[9];
assign y[23] = y2_4[3] & y2_4[5] & y2_4[9];

assign y[24] = y2_4[0] & y2_4[6] & y2_4[9];
assign y[25] = y2_4[1] & y2_4[6] & y2_4[9];
assign y[26] = y2_4[2] & y2_4[6] & y2_4[9];
assign y[27] = y2_4[3] & y2_4[6] & y2_4[9];

assign y[28] = y2_4[0] & y2_4[7] & y2_4[9];
assign y[29] = y2_4[1] & y2_4[7] & y2_4[9];
assign y[30] = y2_4[2] & y2_4[7] & y2_4[9];
assign y[31] = y2_4[3] & y2_4[7] & y2_4[9];

assign y[32] = y2_4[0] & y2_4[4] & y2_4[10];
assign y[33] = y2_4[1] & y2_4[4] & y2_4[10];
assign y[34] = y2_4[2] & y2_4[4] & y2_4[10];
assign y[35] = y2_4[3] & y2_4[4] & y2_4[10];

assign y[36] = y2_4[0] & y2_4[5] & y2_4[10];
assign y[37] = y2_4[1] & y2_4[5] & y2_4[10];
assign y[38] = y2_4[2] & y2_4[5] & y2_4[10];
assign y[39] = y2_4[3] & y2_4[5] & y2_4[10];

assign y[40] = y2_4[0] & y2_4[6] & y2_4[10];
assign y[41] = y2_4[1] & y2_4[6] & y2_4[10];
assign y[42] = y2_4[2] & y2_4[6] & y2_4[10];
assign y[43] = y2_4[3] & y2_4[6] & y2_4[10];

assign y[44] = y2_4[0] & y2_4[7] & y2_4[10];
assign y[45] = y2_4[1] & y2_4[7] & y2_4[10];
assign y[46] = y2_4[2] & y2_4[7] & y2_4[10];
assign y[47] = y2_4[3] & y2_4[7] & y2_4[10];

assign y[48] = y2_4[0] & y2_4[4] & y2_4[11];
assign y[49] = y2_4[1] & y2_4[4] & y2_4[11];
assign y[50] = y2_4[2] & y2_4[4] & y2_4[11];
assign y[51] = y2_4[3] & y2_4[4] & y2_4[11];

assign y[52] = y2_4[0] & y2_4[5] & y2_4[11];
assign y[53] = y2_4[1] & y2_4[5] & y2_4[11];
assign y[54] = y2_4[2] & y2_4[5] & y2_4[11];
assign y[55] = y2_4[3] & y2_4[5] & y2_4[11];

assign y[56] = y2_4[0] & y2_4[6] & y2_4[11];
assign y[57] = y2_4[1] & y2_4[6] & y2_4[11];
assign y[58] = y2_4[2] & y2_4[6] & y2_4[11];
assign y[59] = y2_4[3] & y2_4[6] & y2_4[11];

assign y[60] = y2_4[0] & y2_4[7] & y2_4[11];
assign y[61] = y2_4[1] & y2_4[7] & y2_4[11];
assign y[62] = y2_4[2] & y2_4[7] & y2_4[11];
assign y[63] = y2_4[3] & y2_4[7] & y2_4[11];
endmodule
